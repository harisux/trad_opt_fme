LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.libreria.ALL;

ENTITY filtro_h IS

PORT(A0	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A1	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A2 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A3 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A4 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A5 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A6 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A7 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  CLK	: IN STD_LOGIC;
	  RST : IN STD_LOGIC;
	  SEL1: IN STD_LOGIC;
	  SEL2: IN STD_LOGIC;
	  O1	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  O2	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  O3	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  O4	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END filtro_h;

--------------------------------------------------
--O1: pixel 1/2
--O2: pixel 1/4
--O3: pixel 3/4
--O4: pixel 1
--------------------------------------------------
ARCHITECTURE arq OF filtro_h is


BEGIN

U0: fir_8 PORT MAP(A0=>A0,A1=>A1,A2=>A2,A3=>A3,A4=>A4,A5=>A5,A6=>A6,A7=>A7,CLK=>CLK,RST=>RST,EN=>SEL1,OP=>O4,O=>O1);
U1: fir_7 PORT MAP(A0=>A0,A1=>A1,A2=>A2,A3=>A3,A4=>A4,A5=>A5,A6=>A6,CLK=>CLK,EN=>SEL2,RST=>RST,O=>O2);
U2: fir_7 PORT MAP(A0=>A7,A1=>A6,A2=>A5,A3=>A4,A4=>A3,A5=>A2,A6=>A1,CLK=>CLK,EN=>SEL2,RST=>RST,O=>O3);

END arq;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY fir_8 IS
PORT(A0	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A1	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A2 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A3 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A4 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A5 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A6 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  A7 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  CLK	: IN STD_LOGIC;
	  RST : IN STD_LOGIC;
	  EN	: IN STD_LOGIC;
	  OP	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  O	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END fir_8;

ARCHITECTURE arq OF fir_8 IS

SIGNAL E10: STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL E11: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL E12: STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL E13: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL E14: UNSIGNED(8 DOWNTO 0);
SIGNAL E15: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL E20: SIGNED(11 DOWNTO 0);
SIGNAL E21: SIGNED(9 DOWNTO 0);
SIGNAL E22: STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL E23: STD_LOGIC_VECTOR(12 DOWNTO 0);
SIGNAL E24: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL E30: SIGNED (12 DOWNTO 0);
SIGNAL E31: SIGNED (14 DOWNTO 0);
SIGNAL E32: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL E40: SIGNED(15 DOWNTO 0);
SIGNAL E41: SIGNED(9 DOWNTO 0);
SIGNAL E42: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL R00: STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL R01: STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL R02: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL R03: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL R04: UNSIGNED (8 DOWNTO 0);
SIGNAL R05: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL R10: SIGNED (11 DOWNTO 0);
SIGNAL R11: SIGNED (9 DOWNTO 0);
SIGNAL R12: STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL R13: STD_LOGIC_VECTOR(12 DOWNTO 0);
SIGNAL R14: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL R20: SIGNED (12 DOWNTO 0);
SIGNAL R21: SIGNED (14 DOWNTO 0);
SIGNAL R22: STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN
-- PRIMERA ETAPA FILTRO
	E10 <= (STD_LOGIC_VECTOR(UNSIGNED('0'&A1)+UNSIGNED('0'&A6))&"00");
	E11 <= STD_LOGIC_VECTOR(UNSIGNED('0'&A2)+UNSIGNED('0'&A5));
	E12 <= (STD_LOGIC_VECTOR(E11)&'0');
	E13 <= STD_LOGIC_VECTOR(UNSIGNED('0'&A0)+UNSIGNED('0'&A7));
	E14 <= UNSIGNED('0'&A4)+UNSIGNED('0'&A3);
	E15 <= A3;
	
-- SEGUNDA ETAPA FILTRO
	E20 <= SIGNED('0'&R00)-SIGNED('0'&R01);
	E21 <= SIGNED('0'&R02) + SIGNED('0'&R03);
	E22 <= (STD_LOGIC_VECTOR(R04)&"00000");
	E23 <= (STD_LOGIC_VECTOR(SIGNED('0'&STD_LOGIC_VECTOR(R04))-SIGNED('0'&STD_LOGIC_VECTOR(R02)))&"000");
	E24 <= R05;
	
-- TERCERA ETAPA FILTRO
	E30 <= SIGNED(R10(11)&STD_LOGIC_VECTOR(R10))-SIGNED('0'&STD_LOGIC_VECTOR(R11));
	E31 <= SIGNED('0'&R12)+SIGNED(R13(12)&R13);
	E32 <= R14;
	
-- CUARTA ETAPA FILTRO
	E40 <= SIGNED(R20(12)&STD_LOGIC_VECTOR(R20))+SIGNED('0'&STD_LOGIC_VECTOR(R21));
	E41 <= E40(15 DOWNTO 6);
	E42 <= R22;

--REDONDEAR 
O <= ("11111111") WHEN (E41 > 255) ELSE
	 (OTHERS => '0') WHEN (E41 < 0)  ELSE
	 STD_LOGIC_VECTOR(E41(7 DOWNTO 0));
	 
OP <= E42;

-- REGISTROS
PROCESS(RST,CLK)

BEGIN
	IF (RST='0') THEN 
		R00<=(OTHERS=>'0');
		R01<=(OTHERS=>'0');
		R02<=(OTHERS=>'0');
		R03<=(OTHERS=>'0');
		R04<=(OTHERS=>'0');
		R05<=(OTHERS=>'0');
		R10<=(OTHERS=>'0');
		R11<=(OTHERS=>'0');
		R12<=(OTHERS=>'0');
		R13<=(OTHERS=>'0');
		R14<=(OTHERS=>'0');
		R20<=(OTHERS=>'0');
		R21<=(OTHERS=>'0');
		R22<=(OTHERS=>'0');
	ELSIF RISING_EDGE(CLK) THEN
		IF(EN='1')THEN
			R00 <= E10;
			R01 <= E12;
			R02 <= E11;
			R03 <= E13;
			R04 <= E14;
			R05 <= E15;
			----------
			R10 <= E20;
			R11 <= E21;
			R12 <= E22;
			R13 <= E23;
			R14 <= E24;
			----------
			R20 <= E30;
			R21 <= E31;
			R22 <= E32;
		END IF;
	END IF;
END PROCESS;

END arq;
